package test_pkg;


//import uvm_pkg.sv
	import uvm_pkg::*;
//include uvm_macros.sv
	`include "uvm_macros.svh"
//`include "tb_defs.sv"
`include "src_xtn.sv"
`include "src_agent_config.sv"
`include "dst_agent_config.sv"
`include "env_config.sv"
`include "src_driver.sv"
`include "src_monitor.sv"
`include "src_seqr.sv"
`include "src_agent.sv"
`include "src_agent_top.sv"
`include "src_seq.sv"


`include "dst_xtn.sv"
`include "dst_monitor.sv"
`include "dst_seqr.sv"
`include "dst_seq.sv"
`include "dst_driver.sv"
`include "dst_agent.sv"
`include "dst_agent_top.sv"
`include "virtual_seqr.sv"
`include "virtual_seq.sv"
`include "scoreboard.sv"

`include "env.sv"
`include "vtest_lib.sv"
endpackage






